package ahb_test_pkg;


	import uvm_pkg::*;
	`include "uvm_macros.svh"
	

	`include "ahb_typedefs.sv"
	`include "ahb_master_config.sv"
	`include "ahb_slave_config.sv"
	`include "ahb_env_config.sv"
	
	
	
	`include "ahb_master_xtn.sv"
	`include "ahb_master_driver.sv"
	`include "ahb_master_monitor.sv"	
	`include "ahb_master_sequencer.sv"
	`include "ahb_master_agent.sv"
	`include "ahb_master_agent_top.sv"
	`include "ahb_master_seqs.sv"
	
	
	

	`include "ahb_slave_xtn.sv"
	`include "ahb_slave_driver.sv"
	`include "ahb_slave_monitor.sv"	
	`include "ahb_slave_sequencer.sv"
	`include "ahb_slave_agent.sv"
	`include "ahb_slave_agent_top.sv"
	`include "ahb_slave_seqs.sv"
	
	`include "ahb_virtual_sequencer.sv"
	`include "ahb_virtual_seqs.sv"
	`include "ahb_coverage.sv"
	`include "ahb_tb.sv"
	`include "ahb_vtest_lib.sv"
	

endpackage